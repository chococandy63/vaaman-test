
// Efinity Top-level template
// Version: 2024.1.163
// Date: 2024-10-13 20:24

// Copyright (C) 2013 - 2024 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as /home/trinity/Downloads/efinity/2024.1/project/test_project/test_project.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  test_project
//     #4)  Insert design content.


module test_project
(

);


endmodule

